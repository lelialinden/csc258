module part3 (SW, LEDR, LEDG);
  input [8:0] SW;
  output [8:0] LEDR;
  output [4:0] LEDG;
  
endmodule
