module part7 (SW, KEY)

endmodule
